// Width of fabric 'addr' buses
typedef 32 Wd_Addr;

typedef Bit #(Wd_Addr) Fabric_Addr;
